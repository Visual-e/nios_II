
module nios_cpu (
	clk_clk,
	port_export);	

	input		clk_clk;
	output	[31:0]	port_export;
endmodule
